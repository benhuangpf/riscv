module Decoder(
  input         clock,
  input         reset,
  input  [31:0] io_inst,
  output        io_bundleCtrl_ctrlJump,
  output        io_bundleCtrl_ctrlBranch,
  output        io_bundleCtrl_ctrlRegWrite,
  output        io_bundleCtrl_ctrlLoad,
  output        io_bundleCtrl_ctrlStore,
  output        io_bundleCtrl_ctrlALUSrc,
  output        io_bundleCtrl_ctrlJAL,
  output [3:0]  io_bundleCtrl_ctrlOP,
  output        io_bundleCtrl_ctrlSigned,
  output [1:0]  io_bundleCtrl_ctrlLSType,
  output [4:0]  io_bundleReg_rs1,
  output [4:0]  io_bundleReg_rs2,
  output [4:0]  io_bundleReg_rd,
  output [31:0] io_imm
);
  wire [19:0] _imm_i_T_2 = io_inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 74:12]
  wire [31:0] imm_i = {_imm_i_T_2,io_inst[31:20]}; // @[Cat.scala 31:58]
  wire [31:0] imm_s = {_imm_i_T_2,io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 31:58]
  wire [31:0] imm_b = {_imm_i_T_2,io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] imm_u = {io_inst[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [11:0] _imm_j_T_2 = io_inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 74:12]
  wire [32:0] imm_j = {_imm_j_T_2,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] imm_shamt = {27'h0,io_inst[24:20]}; // @[Cat.scala 31:58]
  wire  _T_11 = io_inst[6:2] == 5'h19; // @[Decoder.scala 72:33]
  wire  _T_13 = io_inst[6:2] == 5'h0; // @[Decoder.scala 78:38]
  wire  _T_15 = io_inst[14:12] == 3'h4; // @[Decoder.scala 82:39]
  wire  _T_17 = io_inst[14:12] == 3'h5; // @[Decoder.scala 82:70]
  wire  _GEN_0 = io_inst[14:12] == 3'h4 | io_inst[14:12] == 3'h5 ? 1'h0 : 1'h1; // @[Decoder.scala 82:84 83:32]
  wire  _T_22 = io_inst[14:12] == 3'h0; // @[Decoder.scala 85:70]
  wire [1:0] _GEN_1 = _T_15 | io_inst[14:12] == 3'h0 ? 2'h0 : 2'h2; // @[Decoder.scala 85:84 86:32]
  wire  _T_25 = io_inst[14:12] == 3'h1; // @[Decoder.scala 88:39]
  wire  _T_28 = io_inst[14:12] == 3'h1 | _T_17; // @[Decoder.scala 88:52]
  wire [1:0] _GEN_2 = io_inst[14:12] == 3'h1 | _T_17 ? 2'h1 : _GEN_1; // @[Decoder.scala 88:84 89:32]
  wire [3:0] _T_39 = {io_inst[30],io_inst[14:12]}; // @[Cat.scala 31:58]
  wire [3:0] _GEN_3 = 4'hd == _T_39 ? 4'hb : 4'h0; // @[Decoder.scala 106:32 95:60]
  wire [3:0] _GEN_4 = 4'h5 == _T_39 ? 4'h9 : _GEN_3; // @[Decoder.scala 102:32 95:60]
  wire [3:0] _GEN_5 = 4'h1 == _T_39 ? 4'h8 : _GEN_4; // @[Decoder.scala 95:60 98:32]
  wire  _T_44 = 3'h0 == io_inst[14:12]; // @[Decoder.scala 111:42]
  wire  _T_45 = 3'h2 == io_inst[14:12]; // @[Decoder.scala 111:42]
  wire  _T_46 = 3'h3 == io_inst[14:12]; // @[Decoder.scala 111:42]
  wire  _T_47 = 3'h4 == io_inst[14:12]; // @[Decoder.scala 111:42]
  wire  _T_48 = 3'h6 == io_inst[14:12]; // @[Decoder.scala 111:42]
  wire  _T_49 = 3'h7 == io_inst[14:12]; // @[Decoder.scala 111:42]
  wire [3:0] _GEN_6 = 3'h7 == io_inst[14:12] ? 4'h4 : 4'h0; // @[Decoder.scala 111:42 135:32]
  wire [3:0] _GEN_7 = 3'h6 == io_inst[14:12] ? 4'h5 : _GEN_6; // @[Decoder.scala 111:42 131:32]
  wire [3:0] _GEN_8 = 3'h4 == io_inst[14:12] ? 4'h7 : _GEN_7; // @[Decoder.scala 111:42 127:32]
  wire [3:0] _GEN_9 = 3'h3 == io_inst[14:12] ? 4'he : _GEN_8; // @[Decoder.scala 111:42 122:32]
  wire  _GEN_10 = 3'h3 == io_inst[14:12] ? 1'h0 : 1'h1; // @[Decoder.scala 111:42 123:36]
  wire [3:0] _GEN_11 = 3'h2 == io_inst[14:12] ? 4'he : _GEN_9; // @[Decoder.scala 111:42 118:32]
  wire [3:0] _GEN_13 = 3'h0 == io_inst[14:12] ? 4'h1 : _GEN_11; // @[Decoder.scala 111:42 114:32]
  wire  _GEN_14 = 3'h0 == io_inst[14:12] | (3'h2 == io_inst[14:12] | _GEN_10); // @[Decoder.scala 111:42]
  wire [31:0] _GEN_15 = io_inst[6:2] == 5'h4 & _T_28 ? imm_shamt : imm_i; // @[Decoder.scala 93:120 110:21 94:21]
  wire [3:0] _GEN_16 = io_inst[6:2] == 5'h4 & _T_28 ? _GEN_5 : _GEN_13; // @[Decoder.scala 93:120]
  wire  _GEN_17 = io_inst[6:2] == 5'h4 & _T_28 | _GEN_14; // @[Decoder.scala 93:120]
  wire [3:0] _GEN_19 = io_inst[6:2] == 5'h0 ? 4'h1 : _GEN_16; // @[Decoder.scala 78:54 80:24]
  wire [31:0] _GEN_20 = io_inst[6:2] == 5'h0 ? imm_i : _GEN_15; // @[Decoder.scala 78:54 81:21]
  wire  _GEN_21 = io_inst[6:2] == 5'h0 ? _GEN_0 : _GEN_17; // @[Decoder.scala 78:54]
  wire [1:0] _GEN_22 = io_inst[6:2] == 5'h0 ? _GEN_2 : 2'h2; // @[Decoder.scala 78:54]
  wire [3:0] _GEN_24 = io_inst[6:2] == 5'h19 ? 4'h1 : _GEN_19; // @[Decoder.scala 72:49 74:24]
  wire [31:0] _GEN_25 = io_inst[6:2] == 5'h19 ? imm_i : _GEN_20; // @[Decoder.scala 72:49 75:21]
  wire  _GEN_26 = io_inst[6:2] == 5'h19 ? 1'h0 : _T_13; // @[Decoder.scala 72:49]
  wire  _GEN_27 = io_inst[6:2] == 5'h19 | _GEN_21; // @[Decoder.scala 72:49]
  wire [1:0] _GEN_28 = io_inst[6:2] == 5'h19 ? 2'h2 : _GEN_22; // @[Decoder.scala 72:49]
  wire  _T_53 = 3'h1 == io_inst[14:12]; // @[Decoder.scala 146:38]
  wire  _T_55 = 3'h5 == io_inst[14:12]; // @[Decoder.scala 146:38]
  wire [3:0] _GEN_29 = _T_49 ? 4'hf : 4'h0; // @[Decoder.scala 146:38 170:28]
  wire  _GEN_30 = _T_49 ? 1'h0 : 1'h1; // @[Decoder.scala 146:38 171:32]
  wire [3:0] _GEN_31 = _T_48 ? 4'he : _GEN_29; // @[Decoder.scala 146:38 165:28]
  wire  _GEN_32 = _T_48 ? 1'h0 : _GEN_30; // @[Decoder.scala 146:38 166:32]
  wire [3:0] _GEN_33 = 3'h5 == io_inst[14:12] ? 4'hf : _GEN_31; // @[Decoder.scala 146:38 161:28]
  wire [3:0] _GEN_35 = _T_47 ? 4'he : _GEN_33; // @[Decoder.scala 146:38 157:28]
  wire [3:0] _GEN_37 = 3'h1 == io_inst[14:12] ? 4'hd : _GEN_35; // @[Decoder.scala 146:38 153:28]
  wire [3:0] _GEN_39 = _T_44 ? 4'hc : _GEN_37; // @[Decoder.scala 146:38 149:28]
  wire  _GEN_40 = _T_44 | (3'h1 == io_inst[14:12] | (_T_47 | (3'h5 == io_inst[14:12] | _GEN_32))); // @[Decoder.scala 146:38]
  wire [1:0] _GEN_41 = _T_22 ? 2'h0 : 2'h2; // @[Decoder.scala 182:49 183:28]
  wire [1:0] _GEN_42 = _T_25 ? 2'h1 : _GEN_41; // @[Decoder.scala 185:49 186:28]
  wire [1:0] _GEN_43 = io_inst[30] ? 2'h2 : 2'h1; // @[Decoder.scala 194:40 195:32 197:32]
  wire [3:0] _GEN_44 = io_inst[30] ? 4'hb : 4'h9; // @[Decoder.scala 219:40 220:32 222:32]
  wire [3:0] _GEN_47 = _T_55 ? _GEN_44 : _GEN_7; // @[Decoder.scala 191:38]
  wire [3:0] _GEN_48 = _T_47 ? 4'h7 : _GEN_47; // @[Decoder.scala 191:38 215:28]
  wire [3:0] _GEN_49 = _T_46 ? 4'h0 : _GEN_48; // @[Decoder.scala 191:38 211:28]
  wire [3:0] _GEN_50 = _T_45 ? 4'he : _GEN_49; // @[Decoder.scala 191:38 206:28]
  wire [3:0] _GEN_51 = _T_53 ? 4'h8 : _GEN_50; // @[Decoder.scala 191:38 202:28]
  wire [3:0] _GEN_52 = _T_44 ? {{2'd0}, _GEN_43} : _GEN_51; // @[Decoder.scala 191:38]
  wire [3:0] _GEN_53 = 5'hc == io_inst[6:2] ? _GEN_52 : 4'h0; // @[Decoder.scala 51:28]
  wire  _GEN_55 = 5'h8 == io_inst[6:2] ? 1'h0 : 1'h1; // @[Decoder.scala 179:26 51:28]
  wire [3:0] _GEN_56 = 5'h8 == io_inst[6:2] ? 4'h1 : _GEN_53; // @[Decoder.scala 180:20 51:28]
  wire [31:0] _GEN_57 = 5'h8 == io_inst[6:2] ? imm_s : 32'h0; // @[Decoder.scala 181:17 51:28]
  wire [1:0] _GEN_58 = 5'h8 == io_inst[6:2] ? _GEN_42 : 2'h2; // @[Decoder.scala 51:28]
  wire  _GEN_59 = 5'h18 == io_inst[6:2] ? 1'h0 : 5'h8 == io_inst[6:2]; // @[Decoder.scala 142:24 51:28]
  wire  _GEN_61 = 5'h18 == io_inst[6:2] ? 1'h0 : _GEN_55; // @[Decoder.scala 144:26 51:28]
  wire [31:0] _GEN_62 = 5'h18 == io_inst[6:2] ? imm_b : _GEN_57; // @[Decoder.scala 145:17 51:28]
  wire [3:0] _GEN_63 = 5'h18 == io_inst[6:2] ? _GEN_39 : _GEN_56; // @[Decoder.scala 51:28]
  wire  _GEN_64 = 5'h18 == io_inst[6:2] ? _GEN_40 : 1'h1; // @[Decoder.scala 51:28]
  wire [1:0] _GEN_65 = 5'h18 == io_inst[6:2] ? 2'h2 : _GEN_58; // @[Decoder.scala 51:28]
  wire  _GEN_66 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] | _GEN_59; // @[Decoder.scala 51:28 70:24]
  wire [3:0] _GEN_68 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] ? _GEN_24 : _GEN_63; // @[Decoder.scala 51:28]
  wire [31:0] _GEN_69 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] ? _GEN_25 : _GEN_62; // @[Decoder.scala 51:28]
  wire  _GEN_71 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] ? _GEN_27 : _GEN_64; // @[Decoder.scala 51:28]
  wire [1:0] _GEN_72 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] ? _GEN_28 : _GEN_65; // @[Decoder.scala 51:28]
  wire  _GEN_73 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] ? 1'h0 : 5'h18 == io_inst[6:2]; // @[Decoder.scala 51:28]
  wire  _GEN_75 = 5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] ? 1'h0 : _GEN_59; // @[Decoder.scala 51:28]
  wire  _GEN_76 = 5'h1b == io_inst[6:2] | _GEN_66; // @[Decoder.scala 51:28 60:24]
  wire  _GEN_77 = 5'h1b == io_inst[6:2] | (5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2]) & _T_11; // @[Decoder.scala 51:28 61:22]
  wire [3:0] _GEN_78 = 5'h1b == io_inst[6:2] ? 4'h1 : _GEN_68; // @[Decoder.scala 51:28 62:20]
  wire [32:0] _GEN_80 = 5'h1b == io_inst[6:2] ? imm_j : {{1'd0}, _GEN_69}; // @[Decoder.scala 51:28 64:17]
  wire  _GEN_81 = 5'h1b == io_inst[6:2] ? 1'h0 : (5'h19 == io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2])
     & _GEN_26; // @[Decoder.scala 51:28]
  wire [1:0] _GEN_83 = 5'h1b == io_inst[6:2] ? 2'h2 : _GEN_72; // @[Decoder.scala 51:28]
  wire  _GEN_84 = 5'h1b == io_inst[6:2] ? 1'h0 : _GEN_73; // @[Decoder.scala 51:28]
  wire  _GEN_86 = 5'h1b == io_inst[6:2] ? 1'h0 : _GEN_75; // @[Decoder.scala 51:28]
  wire [32:0] _GEN_89 = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? {{1'd0}, imm_u} : _GEN_80; // @[Decoder.scala 51:28 56:17]
  assign io_bundleCtrl_ctrlJump = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 1'h0 : _GEN_77; // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlBranch = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 1'h0 : _GEN_84; // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlRegWrite = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] | (5'h1b == io_inst[6:2] | (5'h19 ==
    io_inst[6:2] | 5'h0 == io_inst[6:2] | 5'h4 == io_inst[6:2] | _GEN_61)); // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlLoad = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 1'h0 : _GEN_81; // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlStore = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 1'h0 : _GEN_86; // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlALUSrc = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] | _GEN_76; // @[Decoder.scala 51:28 54:24]
  assign io_bundleCtrl_ctrlJAL = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 1'h0 : 5'h1b == io_inst[6:2]; // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlOP = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 4'h1 : _GEN_78; // @[Decoder.scala 51:28 55:20]
  assign io_bundleCtrl_ctrlSigned = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] | (5'h1b == io_inst[6:2] | _GEN_71); // @[Decoder.scala 51:28]
  assign io_bundleCtrl_ctrlLSType = 5'hd == io_inst[6:2] | 5'h5 == io_inst[6:2] ? 2'h2 : _GEN_83; // @[Decoder.scala 51:28]
  assign io_bundleReg_rs1 = io_inst[19:15]; // @[Decoder.scala 22:32]
  assign io_bundleReg_rs2 = io_inst[24:20]; // @[Decoder.scala 23:32]
  assign io_bundleReg_rd = io_inst[11:7]; // @[Decoder.scala 24:31]
  assign io_imm = _GEN_89[31:0]; // @[Decoder.scala 248:12]
endmodule
