module Alu(
  input         clock,
  input         reset,
  input         io_bundleAluControl_ctrlALUSrc, // @[src/main/scala/examples/Alu.scala 23:16]
  input         io_bundleAluControl_ctrlJAL, // @[src/main/scala/examples/Alu.scala 23:16]
  input  [3:0]  io_bundleAluControl_ctrlOP, // @[src/main/scala/examples/Alu.scala 23:16]
  input         io_bundleAluControl_ctrlSigned, // @[src/main/scala/examples/Alu.scala 23:16]
  input         io_bundleAluControl_ctrlBranch, // @[src/main/scala/examples/Alu.scala 23:16]
  input  [31:0] io_dataRead1, // @[src/main/scala/examples/Alu.scala 23:16]
  input  [31:0] io_dataRead2, // @[src/main/scala/examples/Alu.scala 23:16]
  input  [31:0] io_imm, // @[src/main/scala/examples/Alu.scala 23:16]
  input  [31:0] io_pc, // @[src/main/scala/examples/Alu.scala 23:16]
  output        io_resultBranch, // @[src/main/scala/examples/Alu.scala 23:16]
  output [31:0] io_resultAlu // @[src/main/scala/examples/Alu.scala 23:16]
);
  wire [31:0] oprand1 = io_bundleAluControl_ctrlJAL ? io_pc : io_dataRead1; // @[src/main/scala/examples/Alu.scala 33:19]
  wire [31:0] oprand2 = io_bundleAluControl_ctrlALUSrc ? io_imm : io_dataRead2; // @[src/main/scala/examples/Alu.scala 34:19]
  wire [32:0] _resultAlu_T = oprand1 + oprand2; // @[src/main/scala/examples/Alu.scala 43:34]
  wire [32:0] _resultAlu_T_1 = oprand1 - oprand2; // @[src/main/scala/examples/Alu.scala 46:34]
  wire [31:0] _resultAlu_T_3 = oprand1 & oprand2; // @[src/main/scala/examples/Alu.scala 49:34]
  wire [31:0] _resultAlu_T_4 = oprand1 | oprand2; // @[src/main/scala/examples/Alu.scala 52:34]
  wire [31:0] _resultAlu_T_5 = oprand1 ^ oprand2; // @[src/main/scala/examples/Alu.scala 55:34]
  wire [62:0] _GEN_1 = {{31'd0}, oprand1}; // @[src/main/scala/examples/Alu.scala 58:34]
  wire [62:0] _resultAlu_T_7 = _GEN_1 << oprand2[4:0]; // @[src/main/scala/examples/Alu.scala 58:34]
  wire [31:0] _resultAlu_T_9 = oprand1 >> oprand2[4:0]; // @[src/main/scala/examples/Alu.scala 61:34]
  wire [31:0] _resultAlu_T_10 = io_bundleAluControl_ctrlJAL ? io_pc : io_dataRead1; // @[src/main/scala/examples/Alu.scala 64:35]
  wire [31:0] _resultAlu_T_13 = $signed(_resultAlu_T_10) >>> oprand2[4:0]; // @[src/main/scala/examples/Alu.scala 64:60]
  wire [31:0] _resultBranch_T_1 = io_bundleAluControl_ctrlALUSrc ? io_imm : io_dataRead2; // @[src/main/scala/examples/Alu.scala 67:56]
  wire [32:0] _resultAlu_T_14 = io_pc + io_imm; // @[src/main/scala/examples/Alu.scala 68:32]
  wire  _GEN_0 = io_bundleAluControl_ctrlSigned ? $signed(_resultAlu_T_10) < $signed(_resultBranch_T_1) : oprand1 <
    oprand2; // @[src/main/scala/examples/Alu.scala 76:54 77:34 79:34]
  wire  _GEN_2 = io_bundleAluControl_ctrlBranch & _GEN_0; // @[src/main/scala/examples/Alu.scala 26:35 75:50]
  wire [32:0] _GEN_3 = io_bundleAluControl_ctrlBranch ? _resultAlu_T_14 : {{32'd0}, _GEN_0}; // @[src/main/scala/examples/Alu.scala 75:50 81:27]
  wire  _GEN_4 = io_bundleAluControl_ctrlSigned ? $signed(_resultAlu_T_10) >= $signed(_resultBranch_T_1) : oprand1 >=
    oprand2; // @[src/main/scala/examples/Alu.scala 91:50 92:30 94:30]
  wire  _GEN_5 = 4'hf == io_bundleAluControl_ctrlOP & _GEN_4; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [32:0] _GEN_6 = 4'hf == io_bundleAluControl_ctrlOP ? _resultAlu_T_14 : 33'h0; // @[src/main/scala/examples/Alu.scala 37:40 96:23 27:32]
  wire  _GEN_7 = 4'he == io_bundleAluControl_ctrlOP ? _GEN_2 : _GEN_5; // @[src/main/scala/examples/Alu.scala 37:40]
  wire [32:0] _GEN_8 = 4'he == io_bundleAluControl_ctrlOP ? _GEN_3 : _GEN_6; // @[src/main/scala/examples/Alu.scala 37:40]
  wire  _GEN_9 = 4'hd == io_bundleAluControl_ctrlOP ? $signed(_resultAlu_T_10) != $signed(_resultBranch_T_1) : _GEN_7; // @[src/main/scala/examples/Alu.scala 37:40 71:26]
  wire [32:0] _GEN_10 = 4'hd == io_bundleAluControl_ctrlOP ? _resultAlu_T_14 : _GEN_8; // @[src/main/scala/examples/Alu.scala 37:40 72:23]
  wire  _GEN_11 = 4'hc == io_bundleAluControl_ctrlOP ? $signed(_resultAlu_T_10) == $signed(_resultBranch_T_1) : _GEN_9; // @[src/main/scala/examples/Alu.scala 37:40 67:26]
  wire [32:0] _GEN_12 = 4'hc == io_bundleAluControl_ctrlOP ? _resultAlu_T_14 : _GEN_10; // @[src/main/scala/examples/Alu.scala 37:40 68:23]
  wire [32:0] _GEN_13 = 4'hb == io_bundleAluControl_ctrlOP ? {{1'd0}, _resultAlu_T_13} : _GEN_12; // @[src/main/scala/examples/Alu.scala 37:40 64:23]
  wire  _GEN_14 = 4'hb == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_11; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [32:0] _GEN_15 = 4'h9 == io_bundleAluControl_ctrlOP ? {{1'd0}, _resultAlu_T_9} : _GEN_13; // @[src/main/scala/examples/Alu.scala 37:40 61:23]
  wire  _GEN_16 = 4'h9 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_14; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_17 = 4'h8 == io_bundleAluControl_ctrlOP ? _resultAlu_T_7 : {{30'd0}, _GEN_15}; // @[src/main/scala/examples/Alu.scala 37:40 58:23]
  wire  _GEN_18 = 4'h8 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_16; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_19 = 4'h7 == io_bundleAluControl_ctrlOP ? {{31'd0}, _resultAlu_T_5} : _GEN_17; // @[src/main/scala/examples/Alu.scala 37:40 55:23]
  wire  _GEN_20 = 4'h7 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_18; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_21 = 4'h5 == io_bundleAluControl_ctrlOP ? {{31'd0}, _resultAlu_T_4} : _GEN_19; // @[src/main/scala/examples/Alu.scala 37:40 52:23]
  wire  _GEN_22 = 4'h5 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_20; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_23 = 4'h4 == io_bundleAluControl_ctrlOP ? {{31'd0}, _resultAlu_T_3} : _GEN_21; // @[src/main/scala/examples/Alu.scala 37:40 49:23]
  wire  _GEN_24 = 4'h4 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_22; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_25 = 4'h2 == io_bundleAluControl_ctrlOP ? {{30'd0}, _resultAlu_T_1} : _GEN_23; // @[src/main/scala/examples/Alu.scala 37:40 46:23]
  wire  _GEN_26 = 4'h2 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_24; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_27 = 4'h1 == io_bundleAluControl_ctrlOP ? {{30'd0}, _resultAlu_T} : _GEN_25; // @[src/main/scala/examples/Alu.scala 37:40 43:23]
  wire  _GEN_28 = 4'h1 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_26; // @[src/main/scala/examples/Alu.scala 26:35 37:40]
  wire [62:0] _GEN_29 = 4'h0 == io_bundleAluControl_ctrlOP ? 63'h0 : _GEN_27; // @[src/main/scala/examples/Alu.scala 37:40 39:23]
  assign io_resultBranch = 4'h0 == io_bundleAluControl_ctrlOP ? 1'h0 : _GEN_28; // @[src/main/scala/examples/Alu.scala 37:40 40:26]
  assign io_resultAlu = _GEN_29[31:0]; // @[src/main/scala/examples/Alu.scala 27:32]
endmodule
